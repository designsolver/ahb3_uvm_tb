import uvm_pkg::*;
`include "uvm_macros.svh"

//defines
`include "test/defines.svh"

//rtl
`include "rtl/ahb_if.sv"

//ahb_master_agent
`include "ahb_master_agent/ahb_master_agent_config.sv"
`include "ahb_master_agent/ahb_master_transaction.sv"
`include "ahb_master_agent/sequences/ahb_master_base_sequence.sv"
`include "ahb_master_agent/sequences/ahb_master_idle_sequence.sv"
`include "ahb_master_agent/sequences/ahb_master_incr_sequence.sv"
`include "ahb_master_agent/sequences/ahb_master_single_sequence.sv"
`include "ahb_master_agent/sequences/ahb_master_undeflen_sequence.sv"
`include "ahb_master_agent/sequences/ahb_master_wrap_sequence.sv"
`include "ahb_master_agent/ahb_master_driver.sv"
`include "ahb_master_agent/ahb_master_monitor.sv"
`include "ahb_master_agent/ahb_master_sequencer.sv"
`include "ahb_master_agent/ahb_master_agent.sv"

//ahb_slave_agent
`include "ahb_slave_agent/ahb_slave_agent_config.sv"
`include "ahb_slave_agent/ahb_slave_transaction.sv"
`include "ahb_slave_agent/sequences/ahb_slave_base_sequence.sv"
`include "ahb_slave_agent/sequences/ahb_slave_error_sequence.sv"
`include "ahb_slave_agent/sequences/ahb_slave_okay_sequence.sv"
`include "ahb_slave_agent/ahb_slave_driver.sv"
`include "ahb_slave_agent/ahb_slave_monitor.sv"
`include "ahb_slave_agent/ahb_slave_sequencer.sv"
`include "ahb_slave_agent/ahb_slave_agent.sv"

//ahb_reset_agent
`include "ahb_reset_agent/ahb_reset_agent_config.sv"
`include "ahb_reset_agent/sequences/ahb_reset_sequence.sv"
`include "ahb_reset_agent/sequences/ahb_reset_slave_sequence.sv"
`include "ahb_reset_agent/sequences/ahb_set_sequence.sv"
`include "ahb_reset_agent/ahb_reset_driver.sv"
`include "ahb_reset_agent/ahb_reset_sequencer.sv"
`include "ahb_reset_agent/ahb_reset_agent.sv"

//ahb_env
`include "env/ahb_env_config.sv"
`include "env/vsequences/ahb_base_vseq.sv"
`include "env/ahb_coverage.sv"
`include "env/ahb_env.sv"

//vseq
`include "ahb_vseq.sv"

//test
`include "test/ahb_base_test.sv"
`include "test/init_vseq_from_test.sv"

//top
`include "top.sv"